
package alu_types;

typedef enum logic[2:0] {
  NONE, ADD, SUB, INC, DEC, AND, OR, NOT
} cmd_t /* verilator public */ ;

endpackage : alu_types
