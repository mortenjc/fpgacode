

module register_file(
  input bit clk,
  output bit[31:0] r0,
  output bit[31:0] r1,
  output bit[31:0] r2,
  output bit[31:0] r3,
  output bit[31:0] r4,
  output bit[31:0] r5,
  output bit[31:0] r6,
  output bit[31:0] r7,
  );


always_comb begin

end // always_comb

always_ff @(posedge clk) begin

end // always_ff

endmodule // registers
